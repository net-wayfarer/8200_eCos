# ====================================================================
#
#      ser_mips_bcm33xx.cdl
#
#      eCos serial Broadcom 33xx reference platform configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msieweke
# Original data:  tmichals, dmoseley
# Contributors:
# Date:           2003-07-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

# ====================================================================
# Portions of this software Copyright (c) 2003-2010 Broadcom Corporation
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_MIPS_BCM33XX {
    display       "MIPS BCM33XX reference platform serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_MIPS_BCM33XX

    requires      CYGPKG_ERROR
    include_dir   cyg/io
#    include_files ; # none _exported_ whatsoever
    description   "
           This package contains the serial device drivers for the
           Broadcom 33xx reference platform."

    compile       -library=libextras.a   bcm33xx_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_mips_bcm33xx.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }


cdl_option CYGPKG_IO_SERIAL_MIPS_POLLED_MODE {
    display       "Broadcom 33xx polled mode serial drivers"
    flavor        bool
    default_value 0
    description   "
        If asserted, this option specifies that the serial device
        drivers for the MIPS  should be polled-mode instead of
        interrupt driven."
}

cdl_component CYGPKG_IO_SERIAL_MIPS_BCM33XX_SERIAL_A {
    display       "Broadcom 33xx serial port driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the UART on the 
        Broadcom 33xx."

    cdl_option CYGDAT_IO_SERIAL_MIPS_BCM33XX_SERIAL_A_NAME {
        display       "Device name for Broadcom 33xx serial port"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name on the Broadcom 33xx."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_BCM33XX_SERIAL_A_BAUD {
        display       "Baud rate for the Broadcom 33xx serial port driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 115200
        description   "
            This option specifies the default baud rate (speed) for the 
            Broadcom 33xx serial port."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_BCM33XX_SERIAL_A_BUFSIZE {
        display       "Buffer size for the Broadcom 33xx serial port driver"
        flavor        data
        legal_values  0 to 8192
        default_value 512
        description   "
            This option specifies the size of the internal buffers used
            for the Broadcom 33xx serial port."
    }
}

cdl_component CYGPKG_IO_SERIAL_MIPS_BCM33XX_SERIAL_B {
    display       "Broadcom 33xx serial port driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for the UART on the 
        Broadcom 33xx."

    cdl_option CYGDAT_IO_SERIAL_MIPS_BCM33XX_SERIAL_B_NAME {
        display       "Device name for Broadcom 33xx serial port"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name on the Broadcom 33xx."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_BCM33XX_SERIAL_B_BAUD {
        display       "Baud rate for the Broadcom 33xx serial port driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 115200
        description   "
            This option specifies the default baud rate (speed) for the 
            Broadcom 33xx serial port."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_BCM33XX_SERIAL_B_BUFSIZE {
        display       "Buffer size for the Broadcom 33xx serial port driver"
        flavor        data
        legal_values  0 to 8192
        default_value 512
        description   "
            This option specifies the size of the internal buffers used
            for the Broadcom 33xx serial port."
    }
}

cdl_component CYGPKG_IO_SERIAL_MIPS_BCM33XX_SERIAL_C {
    display       "Broadcom 33xx serial port driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for the UART on the 
        Broadcom 33xx."

    cdl_option CYGDAT_IO_SERIAL_MIPS_BCM33XX_SERIAL_C_NAME {
        display       "Device name for Broadcom 33xx serial port"
        flavor        data
        default_value {"\"/dev/ser2\""}
        description   "
            This option specifies the device name on the Broadcom 33xx."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_BCM33XX_SERIAL_C_BAUD {
        display       "Baud rate for the Broadcom 33xx serial port driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 115200
        description   "
            This option specifies the default baud rate (speed) for the 
            Broadcom 33xx serial port."
    }

    cdl_option CYGNUM_IO_SERIAL_MIPS_BCM33XX_SERIAL_C_BUFSIZE {
        display       "Buffer size for the Broadcom 33xx serial port driver"
        flavor        data
        legal_values  0 to 8192
        default_value 512
        description   "
            This option specifies the size of the internal buffers used
            for the Broadcom 33xx serial port."
    }
}

    cdl_component CYGPKG_IO_SERIAL_MIPS_BCM33XX_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_MIPS_BCM33XX_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_MIPS_BCM33XX_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }
    cdl_component CYGPKG_IO_SERIAL_MIPS_BCM33XX_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_MIPS_BCM33XX_SERIAL_A

        implements CYGINT_IO_SERIAL_TEST_SKIP_9600
        implements CYGINT_IO_SERIAL_TEST_SKIP_14400
        implements CYGINT_IO_SERIAL_TEST_SKIP_38400
        implements CYGINT_IO_SERIAL_TEST_SKIP_57600
        implements CYGINT_IO_SERIAL_TEST_SKIP_PARITY_EVEN
        implements CYGINT_IO_SERIAL_TEST_SKIP_STOP_2

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_MIPS_BCM33XX_SERIAL_A_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"bcm33xx\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF ser_mips_bcm33xx.cdl
